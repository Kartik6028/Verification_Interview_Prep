class packet
    rand bit [31:0] data[8], src;

    constraint c{
        src > 8;
        src <10;
    }

    const bit [31:0] CONG = 42;
    rand bit[31:0] src;
    rand bit congest;
    rand bit [31:0];
    typedef enum  {something, someother, another} stim_e;

    randc bit [1:0] stim_e;

    constraint c_stim {
        len>0;
        len<1000;
        if (congest) {
            dest inside {[cong-10:cong+10]};
            src == cong; //( equivalence operator not assignemnt like =)
        }
        else {
            src inside {0 , [1:10], [10:1000]};

        }

    }

    constraint c_dist {
        src dist {
            0:=40,
            [1:3]:= 60
        }
        /* 0 :40/220;
           1: 60/220;
           2: 60/220;
           3: 60/220;
        */
        dest dist {
            0 :/ 40,
            [1:3] :/ 60
            }
          /*
            0 : 40/100;
            1: 20/100;
            2:  20/100;
            3:  20/100;
          */      
    }

    constraint order {
        low < med;
        med < high;
    }



    constraint c_ins {
        src inside {[low:high]}, //inclusive
        src  inside arr
    }


// SV supports two implication operators for constraints, -> and if
    constrain c_impl {
        check -> addr = 32'hFF; 
       // if check is true then addr must be true, but if check is false then addr can be true or false
       // equal to  (!check || addr)
       // there's also a fully biderectionally visible operator called <->
    }
    // .constraint_mode (0) will switch off a constraint;

    // use with keyword to add extra in-line constraint on the fly on top of existing ones


endclass


packet p;
p = new();

if (!p.randomize()) `UVM_FATAL ()
else transmit (p);


Can you show me how do you write a SV code and assertion check for the spec
Whenever synchronous RESET is set, READY should go low.
2 clocks after every synchronous RESET release, READY should go high.


module xyz
     (
    input clk;
    input rst;
    output rdy;

);

always@ (posedge clk ) begin
    
    if(rst) begin
        rdy =0;
        count =0;        
    end
    else begin
        count <= count+1;
        if (count==2 ) 
        begin
            rdy <=1;
            count<=0;
        end
    
    end

end
    
endmodule


property chk @ (posedge clk )
 (rst) |-> (rdy ==0)
endproperty

property check2 (@ pseedge clk)
 (!rst) |-> #2 rdy;
endproperty


assert chk;

Can you write a python code to parse a file and change the first line first word as 1, 2nd line 2nd word as 2 and so on.
design a traffic controller , control red-green-yellow, input for walk sign. Cycle through RED GREEN YELLOW, whenever input is walk=1, transition to RED LIGHT.


module traffic_controller(
input clk;
input walk;
input rst;
output red;
output green;
output yellow;
);
bit [1:0] state;next_state;
always @(posedge clk)
if (rst)begin
    state<= 2'b00;
    count <=1'b0;

end

else begin 


case (state) begin

2'b00: begin
    state<= 2'b11;
end

2'b01:   //RED
    begin
        count=count+1;
        if ((count == rthreshold )) begin
                state<= 2'b11;
                flag <=0;
         end
         

    end

2'b10:    // YELLOW
    begin
                count=count+1;
              if (count == ythreshold) begin
                state<= 2'b01;
              end

    end

2'b11:   // GREEN
    count=count+1;
    if (count == gthreshold) begin
        state<= 2'b10;
    end

end
endcase


end

always @ (posedge clk )
begin
    if (walk && !flag) begin
        rthreshold= rthreshold +somevalue;
        flag =1; 
    end
    

end




endmodule 



dual port ram - write port and read port, 
 addr;
 data;
 wen;
 ren;

 wen ren
 0   0
 0   1
 1   0
 1   1  // 

 // sequence
    // wr_seq
            // task body
            start_item()
                waddr
                raddr
                data

            finish_item()

            //

    // rd_seq

    

/// DRIVER

//wr_seq.start ()


seq_item_port.get_next_item()
wen=1
ren=1;

drive (pkt);

item_finish


// FIFO - was cannot have a new wr when the fifo is full.

property  fcheck @posedge clk;
$rose(wen) |-> (!full);
endproperty

assert fcheck;

4 different BANKs -
0 - 0 -3 // 
1   4- 7
2   8 - 11
3   12 -15

parameter SIZE =16;
bit [31:0]addr;
add4 [3:0] -  0000
              0011

              0100
              0111


              1000
              1011

              1100
              1111

constraint b1 {
        addr within {  [ start_addr: start_addr + (size*4) ] }

}

constraint ban {
    start_addr[3:2] = 2'b01;

}
    



// write a function take a 32bit input, returns true if value is one hot


function onehot ()

    count = $countones (input)
    if (count ==1) begin
        return true
    else return false

endfunction


return((in & (in -1) ) == 0)

// array of 8 bit vars, constraint for making sure each of the array element is unique 

rand bit [7:0]arr [10];



constraint arr {
    byte data;
    for (int i =0 ; i< arr.size-1 ; i+=) 
        for (int j =1; j<size-1;j++    )
          if (i!=j)  arr[j] != arr[i];
         

    arr [i+1] > arr [i];
}

calculate fifo depth for 100BYTES of data, in a fifo which has no timing consideration. 2 Diff freq 

Read freq = 50 MHZ 
WR FREQ is 150 MHZ
 [ 
    0: BYTE1 
    1: BYTE2
    2: BYTE3  
    3:
    4:
    5:
  ]


design 2 inputs 1 en and 1 input, its intent is to detect pos edge on the input when en is 1, as soon as en is 0 out goes 0


input a
input en
out 

property x @ (posedge clk )

$rose (a) && (en) |-> out; 
endproperty


a en    out
0  0     0  ->  (out) |-> en && $rose(a) 
0  1     a
1  0      
1  1

property y @ (posedge clk )
$fell(en)|-> (out ==0);
endproperty


arr[10]

[1, 2 ,.   .,.. 9,]
val1=0;
equil_index=0





while (lhs!=rhs) begin
    for (int i= equil_index+1; i< size; i++)
         rhs +=  arr[i] ;

    for (int i = 0 ; i=<equil_index; i++) 
        if (equil_index ==0) lhs= 0;
        else  lhs+= arr[i]
    
    if (lhs==rhs) return equil_index;
    else if (equil_index == size-1) return 0;
    else equil_index++;

end

/*

Requirements

Range constraint

All generated addresses must be within the memory map range 0x8000_0000 to 0x8000_FFFF.

Alignment constraint

The address must be 1 KB (1024-byte) aligned.
(In other words, the lower 10 bits of the address must be 0.)

Bank constraint

The 64 KB memory is divided into 4 banks, each of 16 KB (0x4000 bytes).

Bank 0: 0x8000_0000 – 0x8000_3FFF

Bank 1: 0x8000_4000 – 0x8000_7FFF

Bank 2: 0x8000_8000 – 0x8000_BFFF

Bank 3: 0x8000_C000 – 0x8000_FFFF

You must be able to randomize the address only within a specific bank when a variable rand bit [1:0] bank_sel; is set.
For example, if bank_sel == 2'b10, the address should only be from Bank 2.

*/

class packet extends from uvm_transaction;

rand bit [31:0] addr;
rand bit [1:0] bank_sel;

constraint range {

    addr inside {[32'h8000_0000: 32'h8000_FFFF]};
}

constraint alignment {

    addr % 1024 == 0;
}

constraint bank_sel{
   if (bank_sel == 2'b00) addr  inside {[8000_0000:8000_3FFF]};
   if (bank_sel == 2'b01) addr  inside {[8000_4000:8000_7FFF]};
   if (bank_sel == 2'b10) addr  inside {[8000_8000:8000_BFFF]};
   if (bank_sel == 2'b11) addr  inside {[8000_C000:8000_FFFF]};
}

endclass

/*
Specs

addr is 32-bit, must be in [0x4000_0000 : 0x4000_FFFF].

burst_len ∈ {1,2,4,8,16} (beats). Beat size is 4 bytes.

addr must be aligned to burst_len * 4.

The entire burst must not cross a 4 KB page boundary.

Optional targeting: when bank_sel (2 bits) is set, the first beat must be inside the bank window:

Bank 0: [0x4000_0000 : 0x4000_3FFF]

Bank 1: [0x4000_4000 : 0x4000_7FFF]

Bank 2: [0x4000_8000 : 0x4000_BFFF]

Bank 3: [0x4000_C000 : 0x4000_FFFF]


*/

class transaction extends uvm_sequence_item;
rand bit [31:0] addr;
rand bit [3:0] burst_len;


constraint range {
    addr inside {[32'h4000_0000 : 32'h4000_FFFF]};

}

constraint burst_len {
 

    burst_len = $onehot (burst_len);
    //OR
    burst_len == (!(burst_len && (burst_len -1)));
    //OR
    burst_len inside {[4'd1, 4'd2, 4'd4, 4'd8, 4'd16]};
}

constrain aligment {

    addr % (burst_len * 4) == 0;
}

constraint burst_range {

    addr inside {[addr : addr + (burst_len*4) - 1]}
}
endclass


/*
Q2) Whitelist + Blacklist + Weighted Distribution

Constrain an address to allowed regions with weights, block a repeating reserved window, and enforce cacheline alignment.

Specs

addr must land in the whitelist union:
A: [0x9000_0000 : 0x9000_1FFF]
B: [0x9000_4000 : 0x9000_7FFF]
C: [0x9000_C000 : 0x9000_FFFF]

Weights: A:1, B:3, C:2 (i.e., B most likely).

Alignment: 64B (cacheline).

Blacklist pattern: Every 2 KB block reserves the first 256B.
That is, for addr % 2048, the range [0 : 255] is forbidden.

Optional: when is_streaming==1, consecutive randomizations should prefer monotonically increasing addr (hint: use randc/state or a soft constraint).
*/


rand bit [31:0] addr;
constraint range{
    addr dist {[32'h9000_0000: 32'h9000_1FFF] := 1};
    addr dist {[32'h9000_4000: 32'h9000_7FFF] := 3};
    addr dist {[32'h9000_C000: 32'h9000_FFFF] := 2};
}
constraint alignment {
    addr % 8 ==0;
}
constraint forbid {
    if (!(addr % 2048)) {
        addr[11:0] > 12'h0FF;
    }

}
/*

Q3) Page/Offset Build + Set Index Binding

Generate an address from page_num and page_offset, bind index bits to a set_id, and support a “large-page” mode.

Specs

page_num in [0x1000 : 0x1FFF].

Two modes:

large_page==0: page size = 4 KB → page_offset in [0 : 4095].

large_page==1: page size = 2 MB → page_offset in [0 : 2*1024*1024 - 1].

Construct: addr = {page_num, page_offset} only when 4KB pages.
For 2MB pages, ensure resulting addr still falls in [0xA000_0000 : 0xA1FF_FFFF].

Cache set mapping: set_id (6 bits) must equal the index bits of addr[11:6] (i.e., 64 sets, 64B line).

Alignment: 64B lines → addr[5:0] == 0.

Prohibit wraparound across 1MB boundaries for any increment of +N*64B where N∈[0:7].
*/

rand bit [31:0] addr;
rand bit [15:0] page_num;
rand_bit [15:0]page_offset;
rand_bit [31:0]size;
constraint addr_gen {
   if (!large_page) addr = {page_num,page_offset};
   if (large_page)addr inside  {[0xA000_0000: 0xA1FF_FFFF]};
   addr [5:0]==0;
   page_num inside {[16'h1000:16'h1FFF]};

}

constraint page_offset{
    size = large_page? (2*1024*1024): 4096;
    page_offset inside {[16'd0: size-1]};
}

/*
addr must fall in a valid channel and bank range.

Must be aligned to trans_size.

When two consecutive transactions target the same bank, the second one must have a higher address.

You must be able to target a specific channel when force_ch is set.

Transactions must not cross a bank boundary (stay within 64 KB).
CH0 → [0x0000_0000 : 0x0007_FFFF]

CH1 → [0x0008_0000 : 0x000F_FFFF]
*/

rand bit [31:0] addr; 
rand bit [4:0]trans_size;
rand bit channel;
rand bit [2:0]bank_id;
rand bit force_ch;
rand bit [31:0]prev_addr;
constraint addr_range {
    if (force_ch)addr inside {[32'h0000_0000 : 32'h0007_FFFF]}; // select ch0
    else addr inside {[32'h0008_0000: 32'h000F_FFFF]}; // select CH1
}
constraint trans_size {

    trans_size inside {4,8,16,32};
    addr % trans_size ==0;
}
constraint bank_align {
    addr[15:0] + (trans_size * bank_id) <= 16'hFA00; 

}
constraint consecutive {

    if (addr [18:16] == prev_addr [18:16]) {
        addr > prev_addr;
    }
}


/*  
You’re designing a constrained-random generator for DMA transfer descriptors.

Each descriptor includes:

A source address

A destination address

A transfer size

A mode flag (is_secure) that changes which address range is used
*/

rand bit [31:0] src_addr;
rand bit [31:0] dest_addr;
rand bit [7:0]size;
rand bit is_secure;


constraint addr_range {
    src_addr[3:0] == 'b0;
    dest_addr[3:0] == 'b0;


    if (is_secure) {

        src_addr inside {[32'h5000_0000 :  32'h5000_FFFF]};
        dest_addr inside {[ 32'h5000_0000: 32'h5000_FFFF]};

    }

    else {
        src_addr inside {[ 32'h4000_0000: 32'h4000_FFFF]};
        dest_addr inside {[ 32'h4000_0000: 32'h4000_FFFF]};
    }

}

constraint size_rest{
    soft size inside {64,128};
    size inside {16,32,64,128};
    // OR i am giving both options i guess second one below is better ?
    $onehot (size);
    size [3:0] == 'b0;
}

constraint page_boundary{
    (src_addr[11:0] + size) <=  12'hFFF;
    (dest_addr[11:0] + size) <=  12'hFFF;

} 
constraint relation {
    solve src_addr before dest_addr;
    
    if (is_secure) {  
            dest_addr >= src_addr + 12'h100;
    }
   else {
        dest_addr >= src_addr;
   } 

}

constraint non_secure {
    if (!is_secure) {
        dest_addr [9:0] ==src_addr[9:0] + 12'h200;
    }
}


/*
Requirements

There are 8 descriptors, stored in an array addr_q[8].

Each addr_q[i] is a 32-bit address.

All addresses must:

Fall within [0x8000_0000 : 0x8000_0FFF] (4 KB page).

Be 64-byte aligned.

Be unique (no duplicates).

Additionally:

Addresses must be sorted ascending (addr_q[i] < addr_q[i+1]).

The distance between consecutive entries must be at least 128 B apart.

The last entry must not cross the 4 KB boundary.
*/

randc bit [31:0] addr_q [8];

constraint addr_range {

    foreach (addr_q[i]) {
        addr_q[i] inside {[32'h8000_0000 :  32'h8000_0FFF]};
        addr_q[i] [4:0] == 'b0;
        if (i>0)addr_q[i] >= addr_q[i-1] + 8'h80;
        if (i==8)addr_q  <= 12'h1000; 

    }

}
/*
You are writing a constrained-random generator for a queue of packets that are to be sent over a channel.
Each packet has a unique 8-bit ID and a 16-bit payload length.
You must generate a queue of variable length (1–10 packets).
*/

rand bit [7:0] packet_q[$];
rand bit [15:0]payload_length; 
rand bit [3:0]pq_length; 
rand bit [7:0]packet_id;

constraint packetId {

    unique {packet_id};
}

constraint queue_generator {
    soft pq_length inside {4'd8,4'd10};
    payload_length[2:0] =='0;
    pq_length inside {[4'd1:4'd10]};
    (pq_length * 8) < 12'h200;
    foreach (packet_q[i]) {
        if (i<pq_length) {
            packet_q[i].insert(packet_id);
        }
        if (i>0) {
            packet_q[i]>packet_q[0]; 
        }
    }

}



// COVERAGES //

/*
You’re verifying a DMA that supports bursts of 1, 2, 4, 8, and 16 beats, and each beat is 8 bytes.
The 32-bit addr input must always be 8 B-aligned.
You want coverage to ensure you’ve exercised:

All burst lengths,

All page offset regions within a 4 KB page,

And to cross the two, so you can see if large bursts near the 4 KB boundary are tested.

Write a covergroup that:

Samples on every valid transfer (i.e. iff (valid && ready)).

Creates bins for burst_len values {1,2,4,8,16}.

Creates bins for addr[11:0] such that:

low: [0:1023]

mid: [1024:2047]

high: [2048:3071]

near_boundary: [3072:4095]

Cross the two coverpoints.

Mark the combination (burst_len==16 && addr in [3072:4095]) as illegal (since that burst would cross the page boundary).
*/


covergroup cg iff (valid && ready)
    coverpoint addr[2:0];

    coverpoint burst_len [4:0] {
        bins q1 = {1,2,4,8,16};
    }

    

    coverpoint addr[11:0] {

        bins low [] = {[12'd0:12'd1023]};
        bins mid [] = {[12'd1024:12'd2047]};
        bins high[] = {[12'd2048:12'd2071]};
        bins nb [] = {[12'd2072:12'd4095]};


    }


    cross addr, burst_len {
        illegal_bins = burst_len intersect {16} && addr[11:0] intersect {[3072:4095]};
    };

endgroup
/*
🧠 Q2) AXI Write Transaction Coverage

You are verifying an AXI4 write channel.
Each transaction has the following sampled signals:

addr — 32-bit address

burst_len — number of beats (1 – 16)

burst_type — 2-bit value (00 = FIXED, 01 = INCR, 10 = WRAP)

size — 3-bit beat size (e.g., 3’b010 = 4 B/beat)

valid, ready — handshake

You want to create a covergroup that ensures the following are exercised:

1️⃣ All burst types (FIXED, INCR, WRAP)
2️⃣ All burst lengths {1, 4, 8, 16}
3️⃣ All data sizes {1, 2, 4, 8} bytes per beat
4️⃣ Cross coverage of burst_type × size
5️⃣ Mark the combination WRAP + 8 B/beat as illegal (not supported)
6️⃣ Only sample when valid && ready
7️⃣ Optional bonus: add a coverpoint for addr[11:0] (page offset) with bins
  low, mid, high, near_boundary (like before)
*/

covergroup cg with function sample (bit [31:0] addr, bit btype[1:0], bit [3:0] blength, bit [3:0] bpb, bit valid, bit ready );

TYPE:coverpoint btype iff (valid && ready);
LENGTH:coverpoint blength iff (valid && ready) {
    bins legal = {1,4,8,16};
}
DATA_SIZE:coverpoint bpb iff (valid && ready){
    bins legal = {1,2,4,8}
}
cross btype, bpb iff (valid && ready){
    illegal_bins = binsof(TPYE) intersect {01} && binsof(DATA_SIZE) intersect {8};

}
endgroup